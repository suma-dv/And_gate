mailbox gen2drv = new();
mailbox mon2cov = new();
