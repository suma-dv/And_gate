interface intf_gate();
	bit a;
    bit b;
	bit y;
endinterface	
